netcdf profile-Incomplete-MultiDimensional-MultipleProfiles-H.3.2 {
dimensions:
	profile = 142 ;
	alt = 42 ;
variables:
	float lat(profile) ;
		lat:units = "degrees_north" ;
		lat:long_name = "station latitude" ;
		lat:standard_name = "latitude" ;
	float lon(profile) ;
		lon:units = "degrees_east" ;
		lon:long_name = "station longitude" ;
		lon:standard_name = "longitude" ;
	int profile(profile) ;
		profile:cf_role = "profile_id" ;
	int time(profile) ;
		time:long_name = "time" ;
		time:standard_name = "time" ;
		time:units = "seconds since 1990-01-01 00:00:00" ;
		time:missing_value = -999 ;
	float alt(profile, alt) ;
		alt:units = "m" ;
		alt:standard_name = "altitude" ;
		alt:long_name = "height above mean sea level" ;
		alt:positive = "up" ;
		alt:axis = "Z" ;
		alt:missing_value = -999.9f ;
	float temperature(profile, alt) ;
		temperature:long_name = "Air Temperature" ;
		temperature:units = "Celsius" ;
		temperature:coordinates = "time lat lon alt" ;
		temperature:missing_value = -999.9f ;
	float humidity(profile, alt) ;
		humidity:long_name = "Humidity" ;
		humidity:standard_name = "specific_humidity" ;
		humidity:units = "Percent" ;
		humidity:coordinates = "time lat lon alt" ;
		humidity:missing_value = -999.9f ;
	float wind_speed(profile, alt) ;
		wind_speed:long_name = "Wind Speed" ;
		wind_speed:standard_name = "wind_speed" ;
		wind_speed:units = "m/s" ;
		wind_speed:coordinates = "time lat lon alt" ;
		wind_speed:missing_value = -999.9f ;

// global attributes:
		:Conventions = "CF-1.6" ;
		:featureType = "profile" ;
}
