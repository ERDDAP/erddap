netcdf point-H.1 {
dimensions:
	obs = 100 ;
variables:
	double lat(obs) ;
		lat:units = "degrees_north" ;
		lat:long_name = "latitude of the observation" ;
		lat:standard_name = "latitude" ;
	double lon(obs) ;
		lon:units = "degrees_east" ;
		lon:long_name = "longitude of the observation" ;
		lon:standard_name = "longitude" ;
	double alt(obs) ;
		alt:units = "m" ;
		alt:positive = "up" ;
		alt:axis = "Z" ;
		alt:standard_name = "height" ;
	int time(obs) ;
		time:long_name = "time" ;
		time:standard_name = "time" ;
		time:units = "seconds since 1990-01-01 00:00:00" ;
		time:missing_value = -999 ;
	float temperature(obs) ;
		temperature:long_name = "Water Temperature" ;
		temperature:standard_name = "sea_water_temperature" ;
		temperature:units = "Celsius" ;
		temperature:coordinates = "time lat lon alt" ;
		temperature:missing_value = -999.9f ;
	float humidity(obs) ;
		humidity:long_name = "Humidity" ;
		humidity:standard_name = "specific_humidity" ;
		humidity:units = "Percent" ;
		humidity:coordinates = "time lat lon alt" ;
		humidity:missing_value = -999.9f ;

// global attributes:
		:Conventions = "CF-1.6" ;
		:featureType = "point" ;
}
